parameter Num_inp = 222; //number of the cell_units in one row or column  Num_inp x Num_inp MMU 

parameter number_of_calc = 4; //calculator

parameter data_size = 15;  //data size of module

parameter bridge = 25; // bridge for data science

`define DATA_SIZE  10 //data size  = 20
